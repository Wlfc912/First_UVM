package neuron_pkg;
	import uvm_pkg::*;

	`include "neuron_sequencer.sv"
	`include "neuron_monitor.sv"
	`include "neuron_driver.sv"
	`include "neuron_agent.sv"
	`include "neuron_scoreboard.sv"
	`include "neuron_env.sv"
	`include "neuron_test.sv"
endpackage: neuron_pkg